//*****************************************************************************
// Define.vh.
//
// Change History:
//  VER.   Author         DATE              Change Description
//  1.0    Qiwei Wu       Apr. 18, 2020     Initial Release
//*****************************************************************************

`include "Qwi09RegDef.vh"